package pack_ram;
    `include "Transaction.svh"
    `include "Sequencer.svh"
    `include "Driver.svh"
    `include "Monitor.svh"
    `include "Scoreboard.svh"
    `include "Subscriber.svh"
    `include "Environment.svh"
endpackage