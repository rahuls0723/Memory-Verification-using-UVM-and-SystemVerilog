package pack1;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "Ram_Sequence_item.svh"
    `include "Ram_Sequences.svh"
    `include "Ram_Sequencer.svh"
    `include "Ram_Driver.svh"
    `include "Ram_Monitor.svh"
    `include "Ram_Agent.svh"
    `include "Ram_Scoreboard.svh"
    `include "Ram_Subscriber.svh"
    `include "Ram_Env.svh"
    `include "Ram_Test.svh"
endpackage